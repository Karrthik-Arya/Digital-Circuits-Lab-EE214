library ieee;
use ieee.std_logic_1164.all;
package Gates is
  component INVERTER is
   port (A: in std_logic; Y: out std_logic);
  end component INVERTER;

  component AND_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component AND_2;
  
  component AND_3 is
	port (A,B,C: in std_logic; Y: out std_logic);
  end component AND_3;

  component NAND_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component NAND_2;

  component OR_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component OR_2;
  
  component OR_4 is
   port (A, B, C, D: in std_logic; Y: out std_logic);
  end component OR_4;

  component NOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component NOR_2;

  component XOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component XOR_2;

  component XNOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
  end component XNOR_2;

  component HALF_ADDER is
   port (A, B: in std_logic; S, C: out std_logic);
  end component HALF_ADDER;
  
  component Decoder is
   port (A1, A0, E: in std_logic; Y: out std_logic_vector);
  end component Decoder;
  
  component Decoder_3x8 is
   port (A2, A1, A0, E: in std_logic; Y: out std_logic_vector(7 downto 0));
  end component Decoder_3x8;
  
end package Gates;


library ieee;
use ieee.std_logic_1164.all;
entity INVERTER is
   port (A: in std_logic; Y: out std_logic);
end entity INVERTER;

architecture Equations of INVERTER is
begin
   Y <= not A;
end Equations;
  

library ieee;
use ieee.std_logic_1164.all;
entity AND_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity AND_2;


architecture Equations of AND_2 is
begin
   Y <= A and B;
end Equations;
  
library ieee;
use ieee.std_logic_1164.all;
use work.Gates.all;
entity AND_3 is
   port (A, B, C: in std_logic; Y: out std_logic);
end entity AND_3;

architecture Equations of AND_3 is
	signal s1 : std_logic;
begin
   a1 : AND_2 port map(A=> A, B => B, Y => s1);
	a2 : AND_2 port map (A => s1, B => C, Y=> Y);
end Equations;

library ieee;
use ieee.std_logic_1164.all;
entity NAND_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity NAND_2;

architecture Equations of NAND_2 is
begin
   Y <= not (A and B);
end Equations;
  
library ieee;
use ieee.std_logic_1164.all;
entity OR_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity OR_2;

architecture Equations of OR_2 is
begin
   Y <= A or B;
end Equations;

library ieee;
use ieee.std_logic_1164.all;
use work.Gates.all;
entity OR_4 is
   port (A, B, C, D: in std_logic; Y: out std_logic);
end entity OR_4;

architecture Equations of OR_4 is
signal s1, s2: std_logic;
begin
   o1: OR_2 port map (A=>A ,B =>B, Y=> s1);
	o2: OR_2 port map (A=> C, B=> D, Y=> s2);
	o3: OR_2 port map (A=>s1, B=> s2, Y=> Y);
end Equations;

library ieee;
use ieee.std_logic_1164.all;
entity NOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity NOR_2;

architecture Equations of NOR_2 is
begin
   Y <= not (A or B);
end Equations;
  

library ieee;
use ieee.std_logic_1164.all;
entity XOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity XOR_2;

architecture Equations of XOR_2 is
begin
   Y <= A xor B;
end Equations;
  
library ieee;
use ieee.std_logic_1164.all;
entity XNOR_2 is
   port (A, B: in std_logic; Y: out std_logic);
end entity XNOR_2;

architecture Equations of XNOR_2 is
begin
   Y <= not (A xor B);
end Equations;
  
library ieee;
use ieee.std_logic_1164.all;
entity HALF_ADDER is
   port (A, B: in std_logic; S, C: out std_logic);
end entity HALF_ADDER;

architecture Equations of HALF_ADDER is
begin
   S <= (A xor B);
   C <= (A and B);
end Equations;
  
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.Gates.all;
entity Decoder  is
  port (A1, A0, E: in std_logic; Y: out std_logic_vector(3 downto 0));
end entity Decoder;
architecture Struct of Decoder is
  signal N0, N1: std_logic;
begin
  and3: AND_3 port map(A=>A0, B=> A1, C=> E, Y => Y(3));
  not0: INVERTER port map(A=>A0, Y => N0);
  not1: INVERTER port map(A=>A1, Y=>N1);
  and0: AND_3 port map(A=>N0, B=> N1, C=> E, Y=> Y(0));
  and1: AND_3 port map(A=>A0, B=> N1, C=>E, Y=> Y(1));
  and2: AND_3 port map(A=>A1, B => N0, C=>E, Y=> Y(2));
end Struct;

library ieee;
use ieee.std_logic_1164.all;
library work;
use work.Gates.all;
entity Decoder_3x8  is
  port (A2, A1, A0, E: in std_logic; Y: out std_logic_vector(7 downto 0));
end entity Decoder_3x8;
architecture Struct of Decoder_3x8 is
  signal N, S1, S2: std_logic;
begin
  not1: INVERTER port map(A=>A2, Y=>N);
  and1: AND_2 port map(A=>N, B=>E, Y=> S1);
  and2 : AND_2 port map(A=>A2, B=>E, Y=>S2);
  d1: Decoder port map(A0=>A0, A1=>A1, E=> S1, Y=>Y(3 downto 0));
  d2: Decoder port map(A0=>A0, A1=>A1, E=>S2, Y=>Y(7 downto 4));
end Struct;
